`define MODE 1
//1=CRC8 2=CRC12 4=CRC16 8=CRC16-CCITT
`define COUNT 1000
//the number of transaction